
module clock_gater(
    //--------------------------------------------------------------------------
    // Global signals
    //--------------------------------------------------------------------------
    clk,

    //--------------------------------------------------------------------------
    // Input interface
    //--------------------------------------------------------------------------
    i__enable,

    //--------------------------------------------------------------------------
    // Output interface
    //--------------------------------------------------------------------------
    o__gated_clk
);

//------------------------------------------------------------------------------
// Global signals
//------------------------------------------------------------------------------
input  logic                            clk;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Iuput interface
//------------------------------------------------------------------------------
input  logic                            i__enable;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Output interface
//------------------------------------------------------------------------------
output logic                            o__gated_clk;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Signals
//------------------------------------------------------------------------------
logic                                   w__enable_latched;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Generate gated clock
//------------------------------------------------------------------------------
always_latch
begin
    if(clk == 1'b0)
    begin
        w__enable_latched <= i__enable;
    end
end

always_comb
begin
    o__gated_clk = clk & w__enable_latched;
end
//------------------------------------------------------------------------------

endmodule

